--********************************************************
--
-- Notice : 1.   C_S00_AXI_ADDR_WIDTH + 2 >= BRAM_ADDR_SIZE
--          2.   SDK to read BRAM have delay on send times
--         
--********************************************************

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity myip_BRam_ctrl_v1_0 is
	generic (

		-- Parameters of Axi Slave Bus Interface S00_AXI
		C_S00_AXI_DATA_WIDTH	: integer	:= 32;
		C_S00_AXI_ADDR_WIDTH	: integer	:= 32;
		-- Parameters of BRAM Interface
		BRAM_ADDR_SIZE : integer := 19;
		BRAM_DATA_SIZE : integer := 32
		
	);
	port (
		-- block RAM --- Stand Alone mode , Single Port RAM
		addr : out std_logic_vector(BRAM_ADDR_SIZE-1 downto 0) := (others=>'0');  
		clk : out std_logic;
		din : out std_logic_vector(BRAM_DATA_SIZE-1 downto 0):= (others=>'0');  
		dout : in std_logic_vector(BRAM_DATA_SIZE-1 downto 0):= (others=>'0');  
        en : out std_logic := '1';  
        we : out std_logic_vector(0 downto 0) := "0";  --write mode
        rst_active_low : out std_logic := '1';
        
        
		-- Ports of Axi Slave Bus Interface S00_AXI
		s00_axi_aclk	: in std_logic;
		s00_axi_aresetn	: in std_logic;
		s00_axi_awaddr	: in std_logic_vector(C_S00_AXI_ADDR_WIDTH-1 downto 0);
		s00_axi_awprot	: in std_logic_vector(2 downto 0);
		s00_axi_awvalid	: in std_logic;
		s00_axi_awready	: out std_logic;
		s00_axi_wdata	: in std_logic_vector(C_S00_AXI_DATA_WIDTH-1 downto 0);
		s00_axi_wstrb	: in std_logic_vector((C_S00_AXI_DATA_WIDTH/8)-1 downto 0);
		s00_axi_wvalid	: in std_logic;
		s00_axi_wready	: out std_logic;
		s00_axi_bresp	: out std_logic_vector(1 downto 0);
		s00_axi_bvalid	: out std_logic;
		s00_axi_bready	: in std_logic;
		s00_axi_araddr	: in std_logic_vector(C_S00_AXI_ADDR_WIDTH-1 downto 0);
		s00_axi_arprot	: in std_logic_vector(2 downto 0);
		s00_axi_arvalid	: in std_logic;
		s00_axi_arready	: out std_logic;
		s00_axi_rdata	: out std_logic_vector(C_S00_AXI_DATA_WIDTH-1 downto 0);
		s00_axi_rresp	: out std_logic_vector(1 downto 0);
		s00_axi_rvalid	: out std_logic;
		s00_axi_rready	: in std_logic
	); 
end myip_BRam_ctrl_v1_0;

architecture arch_imp of myip_BRam_ctrl_v1_0 is 

	-- component declaration
	component myip_BRam_ctrl_v1_0_S00_AXI is
		generic (
		C_S_AXI_DATA_WIDTH	: integer	:= 32;
		C_S_AXI_ADDR_WIDTH	: integer	:= 4;
		
		BRAM_ADDR_SIZE : integer;
        BRAM_DATA_SIZE : integer
		);
		port (
        
        bram_addr : out std_logic_vector(BRAM_ADDR_SIZE-1 downto 0) := (others=>'0');  
        bram_din : out std_logic_vector(BRAM_DATA_SIZE-1 downto 0);
        bram_dout : in std_logic_vector(BRAM_DATA_SIZE-1 downto 0);
        bram_en : out std_logic := '1';  
        bram_we : out std_logic_vector(0 downto 0) := "1";  --write mode
        
		S_AXI_ACLK	: in std_logic;
		S_AXI_ARESETN	: in std_logic;
		S_AXI_AWADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		S_AXI_AWPROT	: in std_logic_vector(2 downto 0);
		S_AXI_AWVALID	: in std_logic;
		S_AXI_AWREADY	: out std_logic;
		S_AXI_WDATA	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		S_AXI_WSTRB	: in std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
		S_AXI_WVALID	: in std_logic;
		S_AXI_WREADY	: out std_logic;
		S_AXI_BRESP	: out std_logic_vector(1 downto 0);
		S_AXI_BVALID	: out std_logic;
		S_AXI_BREADY	: in std_logic;
		S_AXI_ARADDR	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		S_AXI_ARPROT	: in std_logic_vector(2 downto 0);
		S_AXI_ARVALID	: in std_logic;
		S_AXI_ARREADY	: out std_logic;
		S_AXI_RDATA	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		S_AXI_RRESP	: out std_logic_vector(1 downto 0);
		S_AXI_RVALID	: out std_logic;
		S_AXI_RREADY	: in std_logic
		);
	end component myip_BRam_ctrl_v1_0_S00_AXI;

begin

-- Instantiation of Axi Bus Interface S00_AXI
myip_BRam_ctrl_v1_0_S00_AXI_inst : myip_BRam_ctrl_v1_0_S00_AXI
	generic map (
		C_S_AXI_DATA_WIDTH	=> C_S00_AXI_DATA_WIDTH,
		C_S_AXI_ADDR_WIDTH	=> C_S00_AXI_ADDR_WIDTH,
		BRAM_ADDR_SIZE => BRAM_ADDR_SIZE,
        BRAM_DATA_SIZE => BRAM_DATA_SIZE
	)
	port map (
	   ----BRam port------------------------------------------------
        bram_addr => addr,
        bram_din => din,
        bram_dout => dout,
        bram_en => en,  
        bram_we => we,
        
		S_AXI_ACLK	=> s00_axi_aclk,
		S_AXI_ARESETN	=> s00_axi_aresetn,
		S_AXI_AWADDR	=> s00_axi_awaddr,
		S_AXI_AWPROT	=> s00_axi_awprot,
		S_AXI_AWVALID	=> s00_axi_awvalid,
		S_AXI_AWREADY	=> s00_axi_awready,
		S_AXI_WDATA	=> s00_axi_wdata,
		S_AXI_WSTRB	=> s00_axi_wstrb,
		S_AXI_WVALID	=> s00_axi_wvalid,
		S_AXI_WREADY	=> s00_axi_wready,
		S_AXI_BRESP	=> s00_axi_bresp,
		S_AXI_BVALID	=> s00_axi_bvalid,
		S_AXI_BREADY	=> s00_axi_bready,
		S_AXI_ARADDR	=> s00_axi_araddr,
		S_AXI_ARPROT	=> s00_axi_arprot,
		S_AXI_ARVALID	=> s00_axi_arvalid,
		S_AXI_ARREADY	=> s00_axi_arready,
		S_AXI_RDATA	=> s00_axi_rdata,
		S_AXI_RRESP	=> s00_axi_rresp,
		S_AXI_RVALID	=> s00_axi_rvalid,
		S_AXI_RREADY	=> s00_axi_rready
	);

-----BRam interconnect---------------------------------------------
    clk <= s00_axi_aclk; --BRam clk
    rst_active_low <= s00_axi_aresetn; --BRam reset

end arch_imp;
